module Decoder_3_8(in, out);
	input [2:0] in;
	output [7:0] out;

	wire A, B, C;

	assign out[0] = ~A & ~B & ~C;
	assign out[1] = ~A & ~B & C;
	assign out[2] = ~A & B & ~C;
	assign out[3] = ~A & B & C;
	assign out[4] = A & ~B & ~C;
	assign out[5] = A & ~B & C;
	assign out[6] = A & B & ~C;
	assign out[7] = A & B & C;

endmodule




//Instead of actually writing this, we wrote a program to write it for us.
//Technology!
module Decoder_7_128(in, out);
	input [6:0] in;
	output [127:0] out;
	
	wire A, B, C, D, E, F, G;

	assign out[0] = ~A & ~B & ~C & ~D & ~E & ~F & ~G;
	assign out[1] = ~A & ~B & ~C & ~D & ~E & ~F & G;
	assign out[2] = ~A & ~B & ~C & ~D & ~E & F & ~G;
	assign out[3] = ~A & ~B & ~C & ~D & ~E & F & G;
	assign out[4] = ~A & ~B & ~C & ~D & E & ~F & ~G;
	assign out[5] = ~A & ~B & ~C & ~D & E & ~F & G;
	assign out[6] = ~A & ~B & ~C & ~D & E & F & ~G;
	assign out[7] = ~A & ~B & ~C & ~D & E & F & G;
	assign out[8] = ~A & ~B & ~C & D & ~E & ~F & ~G;
	assign out[9] = ~A & ~B & ~C & D & ~E & ~F & G;
	assign out[10] = ~A & ~B & ~C & D & ~E & F & ~G;
	assign out[11] = ~A & ~B & ~C & D & ~E & F & G;
	assign out[12] = ~A & ~B & ~C & D & E & ~F & ~G;
	assign out[13] = ~A & ~B & ~C & D & E & ~F & G;
	assign out[14] = ~A & ~B & ~C & D & E & F & ~G;
	assign out[15] = ~A & ~B & ~C & D & E & F & G;
	assign out[16] = ~A & ~B & C & ~D & ~E & ~F & ~G;
	assign out[17] = ~A & ~B & C & ~D & ~E & ~F & G;
	assign out[18] = ~A & ~B & C & ~D & ~E & F & ~G;
	assign out[19] = ~A & ~B & C & ~D & ~E & F & G;
	assign out[20] = ~A & ~B & C & ~D & E & ~F & ~G;
	assign out[21] = ~A & ~B & C & ~D & E & ~F & G;
	assign out[22] = ~A & ~B & C & ~D & E & F & ~G;
	assign out[23] = ~A & ~B & C & ~D & E & F & G;
	assign out[24] = ~A & ~B & C & D & ~E & ~F & ~G;
	assign out[25] = ~A & ~B & C & D & ~E & ~F & G;
	assign out[26] = ~A & ~B & C & D & ~E & F & ~G;
	assign out[27] = ~A & ~B & C & D & ~E & F & G;
	assign out[28] = ~A & ~B & C & D & E & ~F & ~G;
	assign out[29] = ~A & ~B & C & D & E & ~F & G;
	assign out[30] = ~A & ~B & C & D & E & F & ~G;
	assign out[31] = ~A & ~B & C & D & E & F & G;
	assign out[32] = ~A & B & ~C & ~D & ~E & ~F & ~G;
	assign out[33] = ~A & B & ~C & ~D & ~E & ~F & G;
	assign out[34] = ~A & B & ~C & ~D & ~E & F & ~G;
	assign out[35] = ~A & B & ~C & ~D & ~E & F & G;
	assign out[36] = ~A & B & ~C & ~D & E & ~F & ~G;
	assign out[37] = ~A & B & ~C & ~D & E & ~F & G;
	assign out[38] = ~A & B & ~C & ~D & E & F & ~G;
	assign out[39] = ~A & B & ~C & ~D & E & F & G;
	assign out[40] = ~A & B & ~C & D & ~E & ~F & ~G;
	assign out[41] = ~A & B & ~C & D & ~E & ~F & G;
	assign out[42] = ~A & B & ~C & D & ~E & F & ~G;
	assign out[43] = ~A & B & ~C & D & ~E & F & G;
	assign out[44] = ~A & B & ~C & D & E & ~F & ~G;
	assign out[45] = ~A & B & ~C & D & E & ~F & G;
	assign out[46] = ~A & B & ~C & D & E & F & ~G;
	assign out[47] = ~A & B & ~C & D & E & F & G;
	assign out[48] = ~A & B & C & ~D & ~E & ~F & ~G;
	assign out[49] = ~A & B & C & ~D & ~E & ~F & G;
	assign out[50] = ~A & B & C & ~D & ~E & F & ~G;
	assign out[51] = ~A & B & C & ~D & ~E & F & G;
	assign out[52] = ~A & B & C & ~D & E & ~F & ~G;
	assign out[53] = ~A & B & C & ~D & E & ~F & G;
	assign out[54] = ~A & B & C & ~D & E & F & ~G;
	assign out[55] = ~A & B & C & ~D & E & F & G;
	assign out[56] = ~A & B & C & D & ~E & ~F & ~G;
	assign out[57] = ~A & B & C & D & ~E & ~F & G;
	assign out[58] = ~A & B & C & D & ~E & F & ~G;
	assign out[59] = ~A & B & C & D & ~E & F & G;
	assign out[60] = ~A & B & C & D & E & ~F & ~G;
	assign out[61] = ~A & B & C & D & E & ~F & G;
	assign out[62] = ~A & B & C & D & E & F & ~G;
	assign out[63] = ~A & B & C & D & E & F & G;
	assign out[64] = A & ~B & ~C & ~D & ~E & ~F & ~G;
	assign out[65] = A & ~B & ~C & ~D & ~E & ~F & G;
	assign out[66] = A & ~B & ~C & ~D & ~E & F & ~G;
	assign out[67] = A & ~B & ~C & ~D & ~E & F & G;
	assign out[68] = A & ~B & ~C & ~D & E & ~F & ~G;
	assign out[69] = A & ~B & ~C & ~D & E & ~F & G;
	assign out[70] = A & ~B & ~C & ~D & E & F & ~G;
	assign out[71] = A & ~B & ~C & ~D & E & F & G;
	assign out[72] = A & ~B & ~C & D & ~E & ~F & ~G;
	assign out[73] = A & ~B & ~C & D & ~E & ~F & G;
	assign out[74] = A & ~B & ~C & D & ~E & F & ~G;
	assign out[75] = A & ~B & ~C & D & ~E & F & G;
	assign out[76] = A & ~B & ~C & D & E & ~F & ~G;
	assign out[77] = A & ~B & ~C & D & E & ~F & G;
	assign out[78] = A & ~B & ~C & D & E & F & ~G;
	assign out[79] = A & ~B & ~C & D & E & F & G;
	assign out[80] = A & ~B & C & ~D & ~E & ~F & ~G;
	assign out[81] = A & ~B & C & ~D & ~E & ~F & G;
	assign out[82] = A & ~B & C & ~D & ~E & F & ~G;
	assign out[83] = A & ~B & C & ~D & ~E & F & G;
	assign out[84] = A & ~B & C & ~D & E & ~F & ~G;
	assign out[85] = A & ~B & C & ~D & E & ~F & G;
	assign out[86] = A & ~B & C & ~D & E & F & ~G;
	assign out[87] = A & ~B & C & ~D & E & F & G;
	assign out[88] = A & ~B & C & D & ~E & ~F & ~G;
	assign out[89] = A & ~B & C & D & ~E & ~F & G;
	assign out[90] = A & ~B & C & D & ~E & F & ~G;
	assign out[91] = A & ~B & C & D & ~E & F & G;
	assign out[92] = A & ~B & C & D & E & ~F & ~G;
	assign out[93] = A & ~B & C & D & E & ~F & G;
	assign out[94] = A & ~B & C & D & E & F & ~G;
	assign out[95] = A & ~B & C & D & E & F & G;
	assign out[96] = A & B & ~C & ~D & ~E & ~F & ~G;
	assign out[97] = A & B & ~C & ~D & ~E & ~F & G;
	assign out[98] = A & B & ~C & ~D & ~E & F & ~G;
	assign out[99] = A & B & ~C & ~D & ~E & F & G;
	assign out[100] = A & B & ~C & ~D & E & ~F & ~G;
	assign out[101] = A & B & ~C & ~D & E & ~F & G;
	assign out[102] = A & B & ~C & ~D & E & F & ~G;
	assign out[103] = A & B & ~C & ~D & E & F & G;
	assign out[104] = A & B & ~C & D & ~E & ~F & ~G;
	assign out[105] = A & B & ~C & D & ~E & ~F & G;
	assign out[106] = A & B & ~C & D & ~E & F & ~G;
	assign out[107] = A & B & ~C & D & ~E & F & G;
	assign out[108] = A & B & ~C & D & E & ~F & ~G;
	assign out[109] = A & B & ~C & D & E & ~F & G;
	assign out[110] = A & B & ~C & D & E & F & ~G;
	assign out[111] = A & B & ~C & D & E & F & G;
	assign out[112] = A & B & C & ~D & ~E & ~F & ~G;
	assign out[113] = A & B & C & ~D & ~E & ~F & G;
	assign out[114] = A & B & C & ~D & ~E & F & ~G;
	assign out[115] = A & B & C & ~D & ~E & F & G;
	assign out[116] = A & B & C & ~D & E & ~F & ~G;
	assign out[117] = A & B & C & ~D & E & ~F & G;
	assign out[118] = A & B & C & ~D & E & F & ~G;
	assign out[119] = A & B & C & ~D & E & F & G;
	assign out[120] = A & B & C & D & ~E & ~F & ~G;
	assign out[121] = A & B & C & D & ~E & ~F & G;
	assign out[122] = A & B & C & D & ~E & F & ~G;
	assign out[123] = A & B & C & D & ~E & F & G;
	assign out[124] = A & B & C & D & E & ~F & ~G;
	assign out[125] = A & B & C & D & E & ~F & G;
	assign out[126] = A & B & C & D & E & F & ~G;
	assign out[127] = A & B & C & D & E & F & G;
	
endmodule