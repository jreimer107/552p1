/* execute.v
* This module takes the data outputs from the decode stage and computes the
* arithmetic output based on the current opcode. It also evaluates the current
* condition based on the current codes in the FLAG register.
* @input instr is the current instruction.
* @input ALUSrc determines whether to use the second Register data or the
*	immediate in calculations.
* @input imm is the immediate generated by the Decode stage.
* @input RegData1 and RegData2 are the Register Data.
* @output alu_out is the result of the calculation.
* @output cond_true is 1 when the condition given in the instruction matches the
* 	values in the flag register.
*/
module execute(clk, rst, instr, ALUSrc, imm, RegData1, RegData2, alu_out,
		ForwardA, ForwardB, alu_out_MEM, WriteData, NVZ);
	input clk, rst;
	input [15:0] instr, imm, RegData1, RegData2;
	input ALUSrc;
	//Forwarding inputs
	input [1:0] ForwardA, ForwardB;
	input [15:0] alu_out_MEM, WriteData;

	output [15:0] alu_out;
	output [2:0] NVZ;

	wire [15:0] alu_in, ALUA, ALUB;
	wire alu_ovfl;

	assign alu_in = ALUSrc ? imm : RegData2;

	//Forwarding nonsense
	assign ALUA = (ForwardA == 2'b00) ? RegData1 :
				  (ForwardA == 2'b01) ? WriteData :
				  						alu_out_MEM;
	assign ALUB = (ForwardB == 2'b00) ? alu_in :
				  (ForwardB == 2'b01) ? WriteData :
				  						alu_out_MEM;

	ALU alu(.A(ALUA), .B(ALUB), .op(instr[15:12]), .out(alu_out),
		.ovfl(alu_ovfl));

	flag_reg FLAG(.clk(clk), .rst(rst), .opcode(instr[15:12]),
		.alu_ovfl(alu_ovfl), .alu_out(alu_out), .NVZ(NVZ));

endmodule
