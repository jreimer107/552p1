module Decoder_4_16(in, out);
	input [2:0] in;
	output [7:0] out;

	wire A, B, C, D;

	assign out[000] = ~A & ~B & ~C & ~D;
	assign out[001] = ~A & ~B & ~C &  D;
	assign out[002] = ~A & ~B &  C & ~D;
	assign out[003] = ~A & ~B &  C &  D;
	assign out[004] = ~A &  B & ~C & ~D;
	assign out[005] = ~A &  B & ~C &  D;
	assign out[006] = ~A &  B &  C & ~D;
	assign out[007] = ~A &  B &  C &  D;
	assign out[008] =  A & ~B & ~C & ~D;
	assign out[009] =  A & ~B & ~C &  D;
	assign out[010] =  A & ~B &  C & ~D;
	assign out[011] =  A & ~B &  C &  D;
	assign out[012] =  A &  B & ~C & ~D;
	assign out[013] =  A &  B & ~C &  D;
	assign out[014] =  A &  B &  C & ~D;
	assign out[015] =  A &  B &  C &  D;

endmodule




//Instead of actually writing this, we wrote a program to write it for us.
//Technology!
module Decoder_7_128(in, out);
	input [6:0] in;
	output [127:0] out;
	
	wire A, B, C, D, E, F, G;

	assign out[000] = ~A & ~B & ~C & ~D & ~E & ~F & ~G;
	assign out[001] = ~A & ~B & ~C & ~D & ~E & ~F &  G;
	assign out[002] = ~A & ~B & ~C & ~D & ~E &  F & ~G;
	assign out[003] = ~A & ~B & ~C & ~D & ~E &  F &  G;
	assign out[004] = ~A & ~B & ~C & ~D &  E & ~F & ~G;
	assign out[005] = ~A & ~B & ~C & ~D &  E & ~F &  G;
	assign out[006] = ~A & ~B & ~C & ~D &  E &  F & ~G;
	assign out[007] = ~A & ~B & ~C & ~D &  E &  F &  G;
	assign out[008] = ~A & ~B & ~C &  D & ~E & ~F & ~G;
	assign out[009] = ~A & ~B & ~C &  D & ~E & ~F &  G;
	assign out[010] = ~A & ~B & ~C &  D & ~E &  F & ~G;
	assign out[011] = ~A & ~B & ~C &  D & ~E &  F &  G;
	assign out[012] = ~A & ~B & ~C &  D &  E & ~F & ~G;
	assign out[013] = ~A & ~B & ~C &  D &  E & ~F &  G;
	assign out[014] = ~A & ~B & ~C &  D &  E &  F & ~G;
	assign out[015] = ~A & ~B & ~C &  D &  E &  F &  G;
	assign out[016] = ~A & ~B &  C & ~D & ~E & ~F & ~G;
	assign out[017] = ~A & ~B &  C & ~D & ~E & ~F &  G;
	assign out[018] = ~A & ~B &  C & ~D & ~E &  F & ~G;
	assign out[019] = ~A & ~B &  C & ~D & ~E &  F &  G;
	assign out[020] = ~A & ~B &  C & ~D &  E & ~F & ~G;
	assign out[021] = ~A & ~B &  C & ~D &  E & ~F &  G;
	assign out[022] = ~A & ~B &  C & ~D &  E &  F & ~G;
	assign out[023] = ~A & ~B &  C & ~D &  E &  F &  G;
	assign out[024] = ~A & ~B &  C &  D & ~E & ~F & ~G;
	assign out[025] = ~A & ~B &  C &  D & ~E & ~F &  G;
	assign out[026] = ~A & ~B &  C &  D & ~E &  F & ~G;
	assign out[027] = ~A & ~B &  C &  D & ~E &  F &  G;
	assign out[028] = ~A & ~B &  C &  D &  E & ~F & ~G;
	assign out[029] = ~A & ~B &  C &  D &  E & ~F &  G;
	assign out[030] = ~A & ~B &  C &  D &  E &  F & ~G;
	assign out[031] = ~A & ~B &  C &  D &  E &  F &  G;
	assign out[032] = ~A &  B & ~C & ~D & ~E & ~F & ~G;
	assign out[033] = ~A &  B & ~C & ~D & ~E & ~F &  G;
	assign out[034] = ~A &  B & ~C & ~D & ~E &  F & ~G;
	assign out[035] = ~A &  B & ~C & ~D & ~E &  F &  G;
	assign out[036] = ~A &  B & ~C & ~D &  E & ~F & ~G;
	assign out[037] = ~A &  B & ~C & ~D &  E & ~F &  G;
	assign out[038] = ~A &  B & ~C & ~D &  E &  F & ~G;
	assign out[039] = ~A &  B & ~C & ~D &  E &  F &  G;
	assign out[040] = ~A &  B & ~C &  D & ~E & ~F & ~G;
	assign out[041] = ~A &  B & ~C &  D & ~E & ~F &  G;
	assign out[042] = ~A &  B & ~C &  D & ~E &  F & ~G;
	assign out[043] = ~A &  B & ~C &  D & ~E &  F &  G;
	assign out[044] = ~A &  B & ~C &  D &  E & ~F & ~G;
	assign out[045] = ~A &  B & ~C &  D &  E & ~F &  G;
	assign out[046] = ~A &  B & ~C &  D &  E &  F & ~G;
	assign out[047] = ~A &  B & ~C &  D &  E &  F &  G;
	assign out[048] = ~A &  B &  C & ~D & ~E & ~F & ~G;
	assign out[049] = ~A &  B &  C & ~D & ~E & ~F &  G;
	assign out[050] = ~A &  B &  C & ~D & ~E &  F & ~G;
	assign out[051] = ~A &  B &  C & ~D & ~E &  F &  G;
	assign out[052] = ~A &  B &  C & ~D &  E & ~F & ~G;
	assign out[053] = ~A &  B &  C & ~D &  E & ~F &  G;
	assign out[054] = ~A &  B &  C & ~D &  E &  F & ~G;
	assign out[055] = ~A &  B &  C & ~D &  E &  F &  G;
	assign out[056] = ~A &  B &  C &  D & ~E & ~F & ~G;
	assign out[057] = ~A &  B &  C &  D & ~E & ~F &  G;
	assign out[058] = ~A &  B &  C &  D & ~E &  F & ~G;
	assign out[059] = ~A &  B &  C &  D & ~E &  F &  G;
	assign out[060] = ~A &  B &  C &  D &  E & ~F & ~G;
	assign out[061] = ~A &  B &  C &  D &  E & ~F &  G;
	assign out[062] = ~A &  B &  C &  D &  E &  F & ~G;
	assign out[063] = ~A &  B &  C &  D &  E &  F &  G;
	assign out[064] =  A & ~B & ~C & ~D & ~E & ~F & ~G;
	assign out[065] =  A & ~B & ~C & ~D & ~E & ~F &  G;
	assign out[066] =  A & ~B & ~C & ~D & ~E &  F & ~G;
	assign out[067] =  A & ~B & ~C & ~D & ~E &  F &  G;
	assign out[068] =  A & ~B & ~C & ~D &  E & ~F & ~G;
	assign out[069] =  A & ~B & ~C & ~D &  E & ~F &  G;
	assign out[070] =  A & ~B & ~C & ~D &  E &  F & ~G;
	assign out[071] =  A & ~B & ~C & ~D &  E &  F &  G;
	assign out[072] =  A & ~B & ~C &  D & ~E & ~F & ~G;
	assign out[073] =  A & ~B & ~C &  D & ~E & ~F &  G;
	assign out[074] =  A & ~B & ~C &  D & ~E &  F & ~G;
	assign out[075] =  A & ~B & ~C &  D & ~E &  F &  G;
	assign out[076] =  A & ~B & ~C &  D &  E & ~F & ~G;
	assign out[077] =  A & ~B & ~C &  D &  E & ~F &  G;
	assign out[078] =  A & ~B & ~C &  D &  E &  F & ~G;
	assign out[079] =  A & ~B & ~C &  D &  E &  F &  G;
	assign out[080] =  A & ~B &  C & ~D & ~E & ~F & ~G;
	assign out[081] =  A & ~B &  C & ~D & ~E & ~F &  G;
	assign out[082] =  A & ~B &  C & ~D & ~E &  F & ~G;
	assign out[083] =  A & ~B &  C & ~D & ~E &  F &  G;
	assign out[084] =  A & ~B &  C & ~D &  E & ~F & ~G;
	assign out[085] =  A & ~B &  C & ~D &  E & ~F &  G;
	assign out[086] =  A & ~B &  C & ~D &  E &  F & ~G;
	assign out[087] =  A & ~B &  C & ~D &  E &  F &  G;
	assign out[088] =  A & ~B &  C &  D & ~E & ~F & ~G;
	assign out[089] =  A & ~B &  C &  D & ~E & ~F &  G;
	assign out[090] =  A & ~B &  C &  D & ~E &  F & ~G;
	assign out[091] =  A & ~B &  C &  D & ~E &  F &  G;
	assign out[092] =  A & ~B &  C &  D &  E & ~F & ~G;
	assign out[093] =  A & ~B &  C &  D &  E & ~F &  G;
	assign out[094] =  A & ~B &  C &  D &  E &  F & ~G;
	assign out[095] =  A & ~B &  C &  D &  E &  F &  G;
	assign out[096] =  A &  B & ~C & ~D & ~E & ~F & ~G;
	assign out[097] =  A &  B & ~C & ~D & ~E & ~F &  G;
	assign out[098] =  A &  B & ~C & ~D & ~E &  F & ~G;
	assign out[099] =  A &  B & ~C & ~D & ~E &  F &  G;
	assign out[100] =  A &  B & ~C & ~D &  E & ~F & ~G;
	assign out[101] =  A &  B & ~C & ~D &  E & ~F &  G;
	assign out[102] =  A &  B & ~C & ~D &  E &  F & ~G;
	assign out[103] =  A &  B & ~C & ~D &  E &  F &  G;
	assign out[104] =  A &  B & ~C &  D & ~E & ~F & ~G;
	assign out[105] =  A &  B & ~C &  D & ~E & ~F &  G;
	assign out[106] =  A &  B & ~C &  D & ~E &  F & ~G;
	assign out[107] =  A &  B & ~C &  D & ~E &  F &  G;
	assign out[108] =  A &  B & ~C &  D &  E & ~F & ~G;
	assign out[109] =  A &  B & ~C &  D &  E & ~F &  G;
	assign out[110] =  A &  B & ~C &  D &  E &  F & ~G;
	assign out[111] =  A &  B & ~C &  D &  E &  F &  G;
	assign out[112] =  A &  B &  C & ~D & ~E & ~F & ~G;
	assign out[113] =  A &  B &  C & ~D & ~E & ~F &  G;
	assign out[114] =  A &  B &  C & ~D & ~E &  F & ~G;
	assign out[115] =  A &  B &  C & ~D & ~E &  F &  G;
	assign out[116] =  A &  B &  C & ~D &  E & ~F & ~G;
	assign out[117] =  A &  B &  C & ~D &  E & ~F &  G;
	assign out[118] =  A &  B &  C & ~D &  E &  F & ~G;
	assign out[119] =  A &  B &  C & ~D &  E &  F &  G;
	assign out[120] =  A &  B &  C &  D & ~E & ~F & ~G;
	assign out[121] =  A &  B &  C &  D & ~E & ~F &  G;
	assign out[122] =  A &  B &  C &  D & ~E &  F & ~G;
	assign out[123] =  A &  B &  C &  D & ~E &  F &  G;
	assign out[124] =  A &  B &  C &  D &  E & ~F & ~G;
	assign out[125] =  A &  B &  C &  D &  E & ~F &  G;
	assign out[126] =  A &  B &  C &  D &  E &  F & ~G;
	assign out[127] =  A &  B &  C &  D &  E &  F &  G;

	
endmodule